// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// Modified for ECE284 Part 2 Project Requirements
`timescale 1ns/1ps

module core_tb;

parameter bw = 4;
parameter psum_bw = 16;
parameter len_kij = 9;
parameter len_onij = 16;
parameter col = 8;
parameter row = 8;
parameter len_nij = 36;

reg clk = 0;
reg reset = 1;

// Increased width to 35 to include mode bit at MSB
wire [34:0] inst_q; 

reg [1:0]  inst_w_q = 0; 
reg [bw*row-1:0] D_xmem_q = 0;
reg CEN_xmem = 1;
reg WEN_xmem = 1;
reg [10:0] A_xmem = 0;
reg CEN_xmem_q = 1;
reg WEN_xmem_q = 1;
reg [10:0] A_xmem_q = 0;
reg CEN_pmem = 1;
reg WEN_pmem = 1;
reg [10:0] A_pmem = 0;
reg CEN_pmem_q = 1;
reg WEN_pmem_q = 1;
reg [10:0] A_pmem_q = 0;
reg ofifo_rd_q = 0;
reg ififo_wr_q = 0;
reg ififo_rd_q = 0;
reg l0_rd_q = 0;
reg l0_wr_q = 0;
reg execute_q = 0;
reg load_q = 0;
reg acc_q = 0;
reg acc = 0;
reg mode = 0; 
reg mode_q = 0;

reg [1:0]  inst_w; 
reg [bw*row-1:0] D_xmem;
reg [psum_bw*col-1:0] answer;

reg ofifo_rd;
reg ififo_wr;
reg ififo_rd;
reg l0_rd;
reg l0_wr;
reg execute;
reg load;

// --- DYNAMIC FILE LOADING VARIABLES ---
reg [8*60:1] data_dir = "./data_files/";  // Directory variable
reg [8*10:1] prefix;                    // Holds "2b_" or "4b_"
reg [8*128:1] w_file_name;
reg [8*128:1] x_file_name;
reg [8*128:1] acc_file_name;
reg [8*128:1] out_file_name;
// --------------------------------------

wire ofifo_valid;
wire [col*psum_bw-1:0] sfp_out;

integer x_file, x_scan_file ; 
integer w_file, w_scan_file ; 
integer acc_file, acc_scan_file ; 
integer out_file, out_scan_file ; 
integer captured_data; 
integer t, i, j, k, kij;
integer ot_idx, max_ot; 
integer error;
integer loop_count;

// Assign mode bit to MSB (Index 34)
assign inst_q[34]   = mode_q; 
assign inst_q[33]   = acc_q;
assign inst_q[32]   = CEN_pmem_q;
assign inst_q[31]   = WEN_pmem_q;
assign inst_q[30:20] = A_pmem_q;
assign inst_q[19]   = CEN_xmem_q;
assign inst_q[18]   = WEN_xmem_q;
assign inst_q[17:7] = A_xmem_q;
assign inst_q[6]    = ofifo_rd_q;
assign inst_q[5]    = ififo_wr_q;
assign inst_q[4]    = ififo_rd_q;
assign inst_q[3]    = l0_rd_q;
assign inst_q[2]    = l0_wr_q;
assign inst_q[1]    = execute_q; 
assign inst_q[0]    = load_q; 


core #(
    .bw(bw),
    .col(col),
    .row(row)
) core_instance (
    .clk(clk), 
    .inst(inst_q),
    .ofifo_valid(ofifo_valid),
    .D_xmem(D_xmem_q), 
    .sfp_out(sfp_out), 
    .reset(reset)
); 

initial begin 
    inst_w   = 0; 
    D_xmem   = 0;
    CEN_xmem = 1;
    WEN_xmem = 1;
    A_xmem   = 0;
    ofifo_rd = 0;
    ififo_wr = 0;
    ififo_rd = 0;
    l0_rd    = 0;
    l0_wr    = 0;
    execute  = 0;
    load     = 0;
    mode     = 0;

    $dumpfile("core_tb.vcd");
    $dumpvars(0,core_tb);

    $display("###################################################");
    $display("############## STARTING PART 2 CHECK ##############");
    $display("###################################################");

    // --- LOOP TWICE: First for 4b, then for 2b ---
    for (loop_count = 0; loop_count < 2; loop_count = loop_count + 1) begin
        // --- SETUP PHASE ---
        if (loop_count == 0) begin
            $display("### STARTING 4-BIT MODE CHECK (Mode=0) ###");
            mode = 0; max_ot = 1; // 4-bit mode: only 1 output tile (8 channels)
            prefix = "4b_";
        end else begin
            $display("### STARTING 2-BIT MODE CHECK (Mode=1) ###");
            mode = 1; max_ot = 2; // 2-bit mode: 2 output tiles (16 channels)
            prefix = "2b_";
        end

        // --- OUTPUT TILE LOOP ---
        for (ot_idx = 0; ot_idx < max_ot; ot_idx = ot_idx + 1) begin
            
            $display(">>> Processing Output Tile %0d <<<", ot_idx);

            A_pmem = 0;

            // Dynamically construct filenames
            $sformat(x_file_name,   "%0s%0sactivation_tile0.txt", data_dir, prefix);
            $sformat(acc_file_name, "%0s%0sacc.txt", data_dir, prefix);
            
            // Generate Out filename with otile index
            if (loop_count == 0) // 4b mode usually doesn't have otile suffix in your gen, adjust if needed
                $sformat(out_file_name, "%0s%0sout.txt", data_dir, prefix);
            else
                $sformat(out_file_name, "%0s%0sout_otile%0d.txt", data_dir, prefix, ot_idx);

            $display("Loading Activation File: %0s", x_file_name);
            
            x_file = $fopen(x_file_name, "r");
            if (x_file == 0) begin $display("ERROR: Could not open file %0s", x_file_name); $finish; end
            
            // Skip headers
            x_scan_file = $fscanf(x_file,"%s", captured_data);
            x_scan_file = $fscanf(x_file,"%s", captured_data);
            x_scan_file = $fscanf(x_file,"%s", captured_data);

            // Reset Sequence
            #0.5 clk = 1'b0;   reset = 1;
            #0.5 clk = 1'b1;

            for (i=0; i<10 ; i=i+1) begin 
                #0.5 clk = 1'b0;
                #0.5 clk = 1'b1; 
            end

            #0.5 clk = 1'b0;   reset = 0;
            #0.5 clk = 1'b1;

            #0.5 clk = 1'b0;   
            #0.5 clk = 1'b1;

            // Activation to xmem 
            for (t=0; t<len_nij; t=t+1) begin  
                #0.5 clk = 1'b0;
                x_scan_file = $fscanf(x_file, "%32b", D_xmem);
                WEN_xmem = 0;
                CEN_xmem = 0;
                if (t>0) A_xmem = A_xmem + 1;
                #0.5 clk = 1'b1;   
            end
            #0.5 clk = 1'b0;  WEN_xmem = 1;  CEN_xmem = 1; A_xmem = 0;
            #0.5 clk = 1'b1; 

            $fclose(x_file);

            // --- KERNEL LOOP ---
            for (kij=0; kij<9; kij=kij+1) begin  
                
                // Generate Weight Filename dynamically with otile index
                $sformat(w_file_name, "%0s%0sweight_itile0_otile%0d_kij%0d.txt", data_dir, prefix, ot_idx, kij);

                w_file = $fopen(w_file_name, "r");
                if (w_file == 0) begin 
                    $display("ERROR: Could not open file %0s", w_file_name); 
                    $finish; 
                end

                // Skip headers
                w_scan_file = $fscanf(w_file,"%s", captured_data);
                w_scan_file = $fscanf(w_file,"%s", captured_data);
                w_scan_file = $fscanf(w_file,"%s", captured_data);

                // Reset before new kernel load (Weight Stationary logic)
                #0.5 clk = 1'b0;    reset = 1;
                #0.5 clk = 1'b1;

                for (i=0; i<10 ; i=i+1) begin 
                    #0.5 clk = 1'b0;
                    #0.5 clk = 1'b1;
                end

                #0.5 clk = 1'b0;    reset = 0;
                #0.5 clk = 1'b1;

                #0.5 clk = 1'b0;    
                #0.5 clk = 1'b1;   

                // Kernel to xmem (Supports SIMD double load)
                A_xmem = 11'b10000000000;
                for (t=0; t<(mode ? col*2 : col); t=t+1) begin  
                    #0.5 clk = 1'b0;
                    w_scan_file = $fscanf(w_file,"%32b", D_xmem);
                    WEN_xmem = 0;
                    CEN_xmem = 0;
                    if (t>0) A_xmem = A_xmem + 1; 
                    #0.5 clk = 1'b1;  
                end

                #0.5 clk = 1'b0;  WEN_xmem = 1;  CEN_xmem = 1; A_xmem = 0;
                #0.5 clk = 1'b1; 

                // Kernel from xmem to L0
                WEN_xmem = 1;
                CEN_xmem = 0;
                l0_wr = 1;
                l0_rd = 0;
                A_xmem = 11'b10000000000;

                for (i=0; i<(mode ? col*2 : col); i=i+1) begin
                    #0.5 clk = 1'b0; 
                    A_xmem = A_xmem + 1; 
                    #0.5 clk = 1'b1; 
                end

                #0.5 clk = 1'b0;
                l0_wr = 0;
                #0.5 clk = 1'b1;

                // Kernel from L0 to PEs
                #0.5 clk = 1'b0;
                l0_rd = 1;
                #0.5 clk = 1'b1;

                for (i=0; i<(mode ? col*2 : col); i=i+1) begin
                    #0.5 clk = 1'b0;
                    load = 1;
                    #0.5 clk = 1'b1; 
                end

                #0.5 clk = 1'b0;  load = 0; l0_rd = 0;
                #0.5 clk = 1'b1;  
            
                // Activation data from xmem to L0 
                WEN_xmem = 1;
                CEN_xmem = 0;
                l0_wr = 1;
                l0_rd = 0;
                A_xmem = 0;

                for (i=0; i<len_nij; i=i+1) begin
                    #0.5 clk = 1'b0; 
                    A_xmem = A_xmem + 1; 
                    #0.5 clk = 1'b1; 
                end

                #0.5 clk = 1'b0; 
                l0_wr = 0; 
                #0.5 clk = 1'b1;

                // Execution start
                #0.5 clk = 1'b0;
                l0_rd = 1;
                #0.5 clk = 1'b1;

                for (i=0; i<len_nij+row+col; i=i+1) begin
                    #0.5 clk = 1'b0;
                    execute = 1;
                    #0.5 clk = 1'b1; 
                end

                // Stop execution 
                #0.5 clk = 1'b0;  execute = 0; l0_rd = 0;
                #0.5 clk = 1'b1;  

                // OFIFO read and p_mem write
                #0.5 clk = 1'b0; 
                ofifo_rd = 1; 
                #0.5 clk = 1'b1;

                #0.5 clk = 1'b0;
                WEN_pmem = 0;
                CEN_pmem = 0;
                #0.5 clk = 1'b1;

                for (t=0; t<len_nij; t=t+1) begin  
                    #0.5 clk = 1'b0;
                    A_pmem = A_pmem + 1;
                    #0.5 clk = 1'b1;  
                end

                #0.5 clk = 1'b0;  WEN_pmem = 1;  CEN_pmem = 1; ofifo_rd = 0; 
                #0.5 clk = 1'b1; 
                
                $fclose(w_file);
            end  // end of kij loop

            // --- VERIFICATION (Per Output Tile) ---
            acc_file = $fopen(acc_file_name, "r"); 
            out_file = $fopen(out_file_name, "r"); 

            if (acc_file == 0) begin $display("ERROR: Missing %0s", acc_file_name); $finish; end
            if (out_file == 0) begin $display("ERROR: Missing %0s", out_file_name); $finish; end

            error = 0;
            $display("############ Verification Start for Output Tile %0d #############", ot_idx); 

            
            for (i=0; i<len_onij+1; i=i+1) begin 
                #0.5 clk = 1'b0; 
                #0.5 clk = 1'b1; 

                if (i>0) begin
                    out_scan_file = $fscanf(out_file,"%128b", answer); 
                    if (sfp_out == answer) begin
                        $display("Output Tile %0d Data %2d matched!", ot_idx, i);
                    end else begin
                        $display("Output Tile %0d Data %2d ERROR!!", ot_idx, i);
                        $display("sfp_out: %128b", sfp_out);
                        $display("answer : %128b", answer);
                        error = 1;
                    end
                end
            
                #0.5 clk = 1'b0; reset = 1;
                #0.5 clk = 1'b1;  
                #0.5 clk = 1'b0; reset = 0;
                #0.5 clk = 1'b1;  

                for (j=0; j<len_kij+1; j=j+1) begin 
                    #0.5 clk = 1'b0;    
                    if (j<len_kij) begin
                        CEN_pmem = 0;
                        WEN_pmem = 1;
                        acc_scan_file = $fscanf(acc_file,"%11b", A_pmem);
                    end else begin
                        CEN_pmem = 1;
                        WEN_pmem = 1;
                    end
                    if (j>0)  acc = 1;  
                    #0.5 clk = 1'b1;    
                end
                #0.5 clk = 1'b0; acc = 0;
                #0.5 clk = 1'b1; 
            end

            if (error == 0) begin
                $display("############ Output Tile %0d PASSED ##############", ot_idx); 
            end else begin
                $display("############ ERROR DETECTED - STOPPING ##############");
                $finish;
            end

            $fclose(acc_file);
            $fclose(out_file);
        
        end // End of ot_idx loop
    
    end // End of loop_count (Run both modes)

    $display("########### Project Part 2 Completed !! ############"); 
    #100 $finish;
end


always @ (posedge clk) begin
   inst_w_q   <= inst_w; 
   D_xmem_q   <= D_xmem;
   CEN_xmem_q <= CEN_xmem;
   WEN_xmem_q <= WEN_xmem;
   A_pmem_q   <= A_pmem;
   CEN_pmem_q <= CEN_pmem;
   WEN_pmem_q <= WEN_pmem;
   A_xmem_q   <= A_xmem;
   ofifo_rd_q <= ofifo_rd;
   acc_q      <= acc;
   ififo_wr_q <= ififo_wr;
   ififo_rd_q <= ififo_rd;
   l0_rd_q    <= l0_rd;
   l0_wr_q    <= l0_wr ;
   execute_q  <= execute;
   load_q     <= load;
   mode_q     <= mode; 
end

endmodule